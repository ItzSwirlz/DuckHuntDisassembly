																																										  																																																																																																																																																																																																																																																										**********  ****                ******																																																																					                     									         																																																																																																											****																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																	    																																							                                                                                 																																																													   																																												    																																	          					                						      																																																																																																																																																																																																																																																																																																																																											  																																																																																															 																																																																																																																																																												        														            																																																						  																																																																																																								             																																																																																			******************												        																																																																													  													     																																							                       																																															        																																																																																																																																																													                                         																																																																						  																																																																									          																										                       																																										    																																																																																																																																																																																																																**************************************																																																																																																																																																																													      																																																																																																																																																																																																		    ********																																																																															   																									   																																																																																																												                  														  																																																																																																																																							  																																																																																																																																																																																																																																																																																																																																																																																																																																																									       																	     						   																																																            																																																				   												  																                         																											    																											********																																																																								        																																																		           																																																										  																									  																																																																																																																																																																																																																										   																																																																								    								    				  					    																																					    								        							                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                																				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ******************************************  ****                          **************************************************************************************************************************************************************************************************************************************************************************************                     *****************                                                                                                                     





















































  



















*********************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************                                                *************************************************************************                                                                    ..........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                        ..............................................................................................................................................................................................................................................................................................................  ............................................................                                    ...........................................................                                                                  ...............................                                  ......... ...........................................................................................................................................................................................................................................................................               ........................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 .................................                                                                                                               ......................................                                                                 .....................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                    ................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ........        ....                                                                                       ....           ........                .........................                                                                                                   .......................................................................................................................................................................................................................................................................................................................................................   ..............................................................................................................................  NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN..............................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             