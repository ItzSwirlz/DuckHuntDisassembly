																																										  																																																																																																																																																																																																																																																										**********  ****************    ******																																																																																																																																																																																																																						****																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																	    																																							                                                                                 																																																																																																												    																																																																						      																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																								******************																																																																																																																																																																																																																																	        																																																																																																																																																																																																																																																																												  																																																																																																																																	  																																																																																																																																																																																																																																																														**************************************																																																																																																																																																																																																																																																																																																																																																																																					    ********																																																																															   																									   																																																																																																																																											  																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																										     																																																																																																																																																																													    																											    																											********																																																																																																																																		           																																																																																																																																																																																																																																																																																																																																																																																																																																																															    												    																																																																																																																																																																																																																																																																								************    **																																																																																																																																																																																																													  																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																							  **************  **************																																																																																																																  													  			************************************************************************  ********************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************     





















































  



















************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************............................................................      ...........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................              ...............................                 ......... ..................................................................................................................................................................................................................................................................................................................................                                                                      ........................................................................   .................................                                                                     ..............................................................   ..............................................................................................................................................................................................................................................................................................................   ...........................................................   .....................................................................................................         .......................   ...................................................   .....................   .................................   ...........               ............................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ....................        .......................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................   ..............................................................................................................................  NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN..............................................                                                                                                                                                                                                                                                             