                                                                                                 																																																																																														                                                                                              										**********                          **																																																														   				                     									         																																																																																																       					  **																																																																					                   																																																		   																																																																																																																																																																																																																																																																																																																																																																																																						    																																							                                                                                 																																	                                  															                                                                                                                       																																		                                               																																																																																																																																																																																											  																																																					  																																																																																				                                                                                                       																																																																						        														            																																																						  																																																																																																								             																																																																																			******************												        																																				   																																						  													     																																							                       																																															        																																																																																																																																																													                                                                                                                                                                                 												          																										                       																																										    																																																																																																																																																																																																																	********************************    **																												     																																																																																																																																												      																																																																																																																																																                  																																		      ******																																																																															   																									   																																    																																							   																																                  								        																																																																																																																																							  																																																																																																																																																																																																																																																																																																																																																																																																																																																									       																	     						   																																																            																																																				   												  																                         																											    																											********																																																																								        	                  																															           																																																										  																									  																																																																																																																																																																																																																										   																																																																								    								    				  					            															  													    								          					                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                																				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ******************************************  ****                          **************************************************************************************************************************************************************************************************************************************************************************************                     *****************                                                                                                                     





















































  



















*********************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************                                                *************************************************************************                                                                    ..........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ............................................................                                    ...........................................................                                                                                                                                                          ...............................                                         ......... ...........................................................................................................................................................................................................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    .................................                                                                                                                              ......................................                                                                 ......................................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ...............   ........................   ...                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ........        ....                                                                                                ....           ........                                                                                                                                                                                                                        ....................................................................................................................................................................................                                                                                                                                                                                       .............................................................................................................  NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN..............................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               