																																										  																																																																																																																																																																																																																																																										**********  ****************    ******																																																																																																																																																																																																																						****																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																	    																																																																													        		                                																																																																																																													    																																																																						      																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																								******************																																																																																																																																																																																																																																	        																																																																																																																																																																																																																																																																												  																																																																																																																																	  																																																																																																																																																																																																																																																														**************************************																																																																																																																																																																																																																																																																																																																																																																																					    ********																																																																															   																									   																																																																																																																																											  																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																										     																																																																																																																																																																													    																											    																											********																																																																																																																																		           																																																																																																																																																																																																																																																																																																																																																																																																																																																															    												    																																																																																																																																																																																																																																																																								************    **																																																																																																																																																																																																													  																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																							  **************  **************																																																																																																																  													  			************************************************************************  ********************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************     





















































  



















************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************............................................................      ...........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................              ...............................                 ......... ..................................................................................................................................................................................................................................................................................................................................                                                                      ........................................................................   .................................                                                                     ..............................................................   ..............................................................................................................................................................................................................................................................................................................   ...........................................................   .....................................................................................................         .......................   ...................................................   .....................   .................................   ...........               ............................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ....................        .......................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................   ..............................................................................................................................  NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN..............................................                                                                                                                                                                                                                                                             