																																										  																																																																																																																																																																																																																																																										**********  ****************    ******																																																																																																																																																																																																																						****																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																	    																																																																													        		                                																																																																																																													    																																																																						      																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																								******************																																																																																																																																																																																																																																	        																																																																																																																																																																																																																																																																												  																																																																																																																																	  																																																																																																																																																																																																																																																														**************************************																																																																																																																																																																																																																																																																																																																																																																																					    ********																																																																															   																									   																																																																																																																																											  																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																										     																																																																																																																																																																													    																											    																											********																																																																																																																																		           																																																																																																																																																																																																																																																																																																																																																																																																																																																															    												    																																																																																																																																																																																																																																																																								************    **																																																																																																																																																																																																													  																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																																							  **************  **************																																																																																																																  													  			************************************************************************  ********************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************     





















































  



















************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************************............................................................      ...........................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................              ...............................      ......... ..................................................................................................................................................................................................................................................................................................................................                                                                      ........................................................................   .................................                                                                     ..............................................................   ..............................................................................................................................................................................................................................................................................................................   .........................................................................................................................................................................   .......................   ...................................................   .....................   .................................   .......................   ............................................................................                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ....................        .......................................................................................................................................................................................................................................................................................................................................................................................................................................................................................................   ..............................................................................................................................  NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN..............................................                                                                                                                                                                                                                                                             